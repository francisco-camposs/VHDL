LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADORSUBTRATOR IS
PORT(

	A,B : IN STD_LOGIC_VECTOR(0 TO 7);
	OP : IN STD_LOGIC;
	S: OUT STD_LOGIC_VECTOR(0 TO 7);
	LUZ1 : OUT STD_LOGIC;
	LUZ2 : OUT STD_LOGIC
	
);
END SOMADORSUBTRATOR;

ARCHITECTURE LOGICA OF SOMADORSUBTRATOR IS
	COMPONENT SOMADORCOMPLETO IS
	PORT(
		Ai, Bi, CARRY_ENTRADA : IN STD_LOGIC;
		S : OUT STD_LOGIC;
		CARRY_SAIDA : OUT STD_LOGIC
	);
	END COMPONENT SOMADORCOMPLETO;
	
	COMPONENT DECODIFICADOR1X2 IS
	PORT (
		A : IN STD_LOGIC;
		S1, S2 : OUT STD_LOGIC
	); 
	END COMPONENT DECODIFICADOR1X2;
	
	SIGNAL INVERSOR: STD_LOGIC_VECTOR(0 TO 7);
	SIGNAL CARRY: STD_LOGIC_VECTOR(0 TO 7);
	
BEGIN

	INVERSOR(0) <= OP XOR B(0);
	G1 : SOMADORCOMPLETO PORT MAP (A(0),B(0),OP, S(0), CARRY(0));
	
	INVERSOR(1) <= OP XOR B(1);
	G2 : SOMADORCOMPLETO PORT MAP (A(1),B(1),CARRY(0), S(1), CARRY(1));
	
	INVERSOR(2) <= OP XOR B(2);
	G3 : SOMADORCOMPLETO PORT MAP (A(2),B(2),CARRY(1), S(2), CARRY(2));
	
	INVERSOR(3) <= OP XOR B(3);
	G4 : SOMADORCOMPLETO PORT MAP (A(3),B(3),CARRY(2), S(3), CARRY(3));
	
	INVERSOR(4) <= OP XOR B(4);
	G5 : SOMADORCOMPLETO PORT MAP (A(4),B(4),CARRY(3), S(4), CARRY(4));
	
	INVERSOR(5) <= OP XOR B(5);
	G6 : SOMADORCOMPLETO PORT MAP (A(5),B(5),CARRY(4), S(5), CARRY(5));
	
	INVERSOR(6) <= OP XOR B(6);
	G7 : SOMADORCOMPLETO PORT MAP (A(6),B(6),CARRY(5), S(6), CARRY(6));
	
	INVERSOR(7) <= OP XOR B(7);
	G8 : SOMADORCOMPLETO PORT MAP (A(7),B(7),CARRY(6), S(7), CARRY(7));
	
	G9 : DECODIFICADOR1X2 PORT MAP (OP, LUZ1, LUZ2);


END LOGICA;