LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODIFICADOR1X2 IS
PORT (
	A: IN STD_LOGIC;
	S1, S2 : OUT STD_LOGIC
);
END DECODIFICADOR1X2;

ARCHITECTURE LOGICA OF DECODIFICADOR1X2 IS
BEGIN

	S1 <= NOT(A);
	S2 <= A;

END;