LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY A_NAND_B IS
PORT (
	a, b : IN STD_LOGIC;
	x : OUT STD_LOGIC
);
END A_NAND_B;

ARCHITECTURE LOGICA1 OF A_NAND_B IS
BEGIN
	X <= NOT(A AND B);
END LOGICA1;