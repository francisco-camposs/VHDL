LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY A_OR_B IS
PORT (
	a, b : IN STD_LOGIC;
	x : OUT STD_LOGIC
);
END A_OR_B;

ARCHITECTURE LOGICA2 OF A_OR_B IS
BEGIN
	X <= A OR B;
END LOGICA2;