LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PrimeiraColuna IS
PORT(
	A1, B1 : IN STD_LOGIC;
	S1 : OUT STD_LOGIC;
	C1 : OUT STD_LOGIC
);
END PrimeiraColuna;

ARCHITECTURE LOGICA OF PrimeiraColuna IS
BEGIN
	S1 <= A1 XOR B1;
	C1 <= A1 AND B1;
END LOGICA;