LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUBTRATOR IS 
PORT (
	A1, A2 : IN STD_LOGIC_VECTOR(0 TO 3);
	S1 : OUT STD_LOGIC_VECTOR(0 TO 3);
	OVERFLOW : OUT STD_LOGIC
);
END SUBTRATOR;

ARCHITECTURE Aula10Exercicio1 of SUBTRATOR is

COMPONENT SOMADOR4BITS
PORT(
	A1,A2 : IN STD_LOGIC_VECTOR(0 TO 3);
	S1: OUT STD_LOGIC_VECTOR(0 TO 3);
	OVERFLOW_SUBTRACAO : OUT STD_LOGIC;
	OVERFLOW : OUT STD_LOGIC
);
END COMPONENT;

SIGNAL AUX0 : STD_LOGIC_VECTOR(0 TO 3);
SIGNAL AUX1 : STD_LOGIC_VECTOR(0 TO 3);
SIGNAL AUX2 : STD_LOGIC_VECTOR(0 TO 3);

BEGIN

	P1 : SOMADOR4BITS PORT MAP ("0001", "0001", S1,AUX0(0), AUX0(1));
	

END Aula10Exercicio1;




