LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NXOR IS
PORT (
	A, B, CARRY : IN STD_LOGIC;
	S : OUT STD_LOGIC
);
END NXOR;

ARCHITECTURE LOGICA OF NXOR IS
BEGIN

S <= (A AND NOT(B) AND NOT(CARRY)) OR (NOT(A) AND NOT(B) AND CARRY) OR (A AND B AND CARRY) OR (NOT(A) AND B AND NOT(CARRY));

END LOGICA;