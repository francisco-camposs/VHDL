LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Aula4Exercicio1 IS
PORT (
	E1 : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	S1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END Aula4Exercicio1;

ARCHITECTURE AAND OF Aula4Exercicio1 IS
	SUBTYPE BYTE IS  STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL B1 : BYTE := "10011001";
BEGIN
	E1(0) <= B1(0);
	E1(1) <= B1(1);
	E1(2) <= B1(2);
	E1(3) <= B1(3);
	E1(4) <= B1(4);
	E1(5) <= B1(5);
	E1(6) <= B1(6);
	E1(7) <= B1(7);
	
	S1(0) <= E1(0);
	S1(1) <= E1(1);
	S1(2) <= E1(2);
	S1(3) <= E1(3);
	S1(4) <= E1(4);
	S1(5) <= E1(5);
	S1(6) <= E1(6);
	S1(7) <= E1(7);

END AAND;