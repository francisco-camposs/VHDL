LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY A_NOR_B IS
PORT (
	a, b : IN STD_LOGIC;
	x : OUT STD_LOGIC
);
END A_NOR_B;

ARCHITECTURE LOGICA OF A_NOR_B IS
BEGIN
	X <= NOT(A OR B);
END LOGICA;