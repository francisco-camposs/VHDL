LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR4BITS IS
PORT(
	A1, A2 : IN STD_LOGIC_VECTOR(0 TO 3);
	S1 : OUT STD_LOGIC_VECTOR(0 TO 3);
	OVERFLOW_SUBTRACAO : OUT STD_LOGIC;
	OVERFLOW : OUT STD_LOGIC
);
END SOMADOR4BITS;

ARCHITECTURE  LOGICA OF SOMADOR4BITS IS

COMPONENT PrimeiraColuna is
PORT(
	A1, B1 : IN STD_LOGIC;
	S1 : OUT STD_LOGIC;
	C1 : OUT STD_LOGIC
);
END COMPONENT;

COMPONENT DemaisColunas is
PORT(
	A1, B1, C0: IN STD_LOGIC;
	S1 : OUT STD_LOGIC;
	C1 : OUT STD_LOGIC
);
END COMPONENT;

SIGNAL SIG0 : STD_LOGIC_VECTOR(0 TO 3);

BEGIN

	P1 : PrimeiraColuna PORT MAP (A1(0), A2(0), S1(0), SIG0(0));
	P2 : DemaisColunas PORT MAP (A1(1), A2(1), SIG0(0) , S1(1), SIG0(1));
	P3 : DemaisColunas PORT MAP (A1(2), A2(2), SIG0(1) , S1(2), SIG0(2));
	P4 : DemaisColunas PORT MAP (A1(3), A2(3), SIG0(2), S1(3), SIG0(3));
	OVERFLOW_SUBTRACAO <= SIG0(2);
	OVERFLOW <= SIG0(3);

END;