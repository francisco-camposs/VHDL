LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUBTRATOR IS 
PORT (
	A1, A2 : IN STD_LOGIC_VECTOR(0 TO 3);
	TESTE : IN STD_LOGIC;
	S1 : OUT STD_LOGIC_VECTOR(0 TO 3);
	OVERFLOW : OUT STD_LOGIC
);
END SUBTRATOR;

ARCHITECTURE Aula10Exercicio1 of SUBTRATOR is

COMPONENT SOMADORCOMPLETO IS
PORT(
	Ai, Bi, CARRY_ENTRADA : IN STD_LOGIC;
	S : OUT STD_LOGIC;
	CARRY_SAIDA : OUT STD_LOGIC
);
END COMPONENT SOMADORCOMPLETO;

SIGNAL CARRY1 : STD_LOGIC;
SIGNAL CARRY2 : STD_LOGIC;
SIGNAL CARRY3 : STD_LOGIC;
SIGNAL CARRY4 : STD_LOGIC;


BEGIN

	G1 : SOMADORCOMPLETO PORT MAP (A1(0), NOT(A2(0)), '1', S1(0), CARRY1);
	G2 : SOMADORCOMPLETO PORT MAP (A1(1), NOT(A2(1)), CARRY1, S1(1), CARRY2);
	G3 : SOMADORCOMPLETO PORT MAP (A1(2), NOT(A2(2)), CARRY2, S1(2), CARRY3);
	G4 : SOMADORCOMPLETO PORT MAP (A1(3), NOT(A2(3)), CARRY3, S1(3), CARRY4);
	OVERFLOW <= NOT((NOT(CARRY3) AND NOT (CARRY3)) OR (CARRY4 AND CARRY3));

END Aula10Exercicio1;
