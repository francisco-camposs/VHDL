LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY DemaisColunas is
PORT(
	A1, B1, C0: IN STD_LOGIC;
	S1 : OUT STD_LOGIC;
	C1 : OUT STD_LOGIC
);
END DemaisColunas;

ARCHITECTURE LOGICA OF DemaisColunas IS
BEGIN

	S1 <= A1 XOR B1 XOR C0;
	C1 <= (A1 AND B1) OR (C0 AND (B1 XOR A1));

END LOGICA;