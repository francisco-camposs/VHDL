LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NOT_A IS
PORT (
	a: IN STD_LOGIC;
	x : OUT STD_LOGIC
);
END NOT_A;

ARCHITECTURE LOGICA2 OF NOT_A IS
BEGIN
	X <= NOT A;
END LOGICA2;