LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Aula4Exercicio1 IS 
PORT (
	A1 : IN BIT_VECTOR(3 DOWNTO 0);
	B1 : OUT BIT_VECTOR(3 DOWNTO 0)
);
END Aula4Exercicio1;

ARCHITECTURE USAR OF Aula4Exercicio1 IS
	SUBTYPE BARRAMENTO IS BIT_VECTOR(3 DOWNTO 0);
	SIGNAL BARRA : BARRAMENTO;
BEGIN

	BARRA(0) <= A1(0);
	BARRA(1) <= A1(1);
	BARRA(2) <= A1(2);
	BARRA(3) <= A1(3);
	B1(0) <=  BARRA(0);
	B1(1) <=  BARRA(1);
	B1(2) <=  BARRA(2);
	B1(3) <=  BARRA(3);

END USAR;