LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SomadorCompleto IS
PORT (
	Ai, Bi, CARRY_ENTRADA : IN STD_LOGIC;
	S : OUT STD_LOGIC;
	CARRY_SAIDA : out STD_LOGIC
);
END SomadorCompleto;

ARCHITECTURE LOGICA OF SOMADORCOMPLETO IS
	
	COMPONENT NXOR IS
	PORT (
		A, B, CARRY : IN STD_LOGIC;
		S : OUT STD_LOGIC
	);
	END COMPONENT NXOR;

BEGIN

	G1: NXOR PORT MAP (Ai, Bi, CARRY_ENTRADA, S);
	CARRY_SAIDA <= (Bi and CARRY_ENTRADA) or (Ai and CARRY_ENTRADA) or (Ai and Bi);

END LOGICA;