LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPARADOR1BIT IS
	PORT ( 
	A, B : IN STD_LOGIC;
	X, Y, Z : OUT STD_LOGIC );
END COMPARADOR1BIT;

ARCHITECTURE LOGICA OF COMPARADOR1BIT IS
BEGIN
	X <= A XNOR B;
	Y <= A AND (NOT B);
	Z <= (NOT A) AND B;
END LOGICA;