LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EXERCICIO2 IS
PORT (
	A,B,C : IN STD_LOGIC_VECTOR(0 TO 7);
	S : OUT STD_LOGIC_VECTOR(0 TO 7)
);
END EXERCICIO2;

ARCHITECTURE LOGICA OF EXERCICIO2 IS
BEGIN

	S(0 TO 7) <= A(0 TO 7) xnor B(0 TO 7);

END LOGICA;