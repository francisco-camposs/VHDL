LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY circuito IS
PORT (
	a, b, c, d: IN STD_LOGIC;
	x: OUT STD_LOGIC
);
END circuito;

ARCHITECTURE ESTRUTURAL OF CIRCUITO IS
	COMPONENT A_AND_B IS
	PORT (
		A,B : IN STD_LOGIC;
		X : OUT STD_LOGIC
	);
	END COMPONENT A_AND_B;
	
	COMPONENT A_OR_B IS
	PORT (
		A, B : IN STD_LOGIC;
		X : OUT STD_LOGIC
	);
	END COMPONENT A_OR_B;
	
	COMPONENT A_NOR_B IS
	PORT (
		A, B : IN STD_LOGIC;
		X : OUT STD_LOGIC
	);
	END COMPONENT A_NOR_B;
	
	COMPONENT A_NAND_B IS
	PORT (
		A, B : IN STD_LOGIC;
		X : OUT STD_LOGIC
	);
	END COMPONENT A_NAND_B;
	
	COMPONENT NOT_A IS
	PORT (
		A: IN STD_LOGIC;
		X : OUT STD_LOGIC
	);
	END COMPONENT NOT_A;
	
	SIGNAL AUX1 : STD_LOGIC;
	SIGNAL AUX2 : STD_LOGIC;
	SIGNAL AUX3 : STD_LOGIC;
	SIGNAL AUX4 : STD_LOGIC;
	SIGNAL AUX5 : STD_LOGIC;
	SIGNAL AUX6 : STD_LOGIC;
	SIGNAL AUX7 : STD_LOGIC;
	SIGNAL AUX8 : STD_LOGIC;
	SIGNAL AUX8_5 : STD_LOGIC;
	SIGNAL AUX9 : STD_LOGIC;


BEGIN

	G1 : A_AND_B PORT MAP (a, b, AUX1);
	G2 : A_NAND_B PORT MAP (b, c, AUX2);
	G3 : NOT_A PORT MAP (B, AUX3);
	G4 : NOT_A PORT MAP (C, AUX4);
	G5 : A_AND_B PORT MAP (AUX3, AUX4, AUX5);
	G6 : A_OR_B PORT MAP (AUX5, C, AUX6);
	G7 : A_OR_B PORT MAP (AUX1, AUX2, AUX7);
	G8 : NOT_A PORT MAP (AUX6, AUX8);
	G8_5 : NOT_A PORT MAP (D, AUX8_5);
	G9 : A_AND_B PORT MAP (AUX8_5, AUX8, AUX9);
	G10 : A_OR_B PORT MAP (AUX7, AUX9, X);
	

END ESTRUTURAL; 
